`ifndef CONST
`define CONST

`define MODE_WIDTH 2
`define LABEL_WIDTH 5
`define HV_DIMENSION 1000
`define DISTANCE_WIDTH 10
`define CLASSES 21
`define INPUT_CHANNELS 64
`define CHANNEL_WIDTH 6
`define RAW_WIDTH 15
`define SPATIAL_WIDTH 13
`define SPATIAL_N 8
`define SPATIAL_DIMENSION `HV_DIMENSION/`SPATIAL_N
`define NGRAM_SIZE 5
`define SBUFFER_DEPTH 32
`define FEATWIN_SIZE 50
`define MAX_BUNDLE_CYCLES 80
`define BUNDLE_NGRAMS_WIDTH 7
`define HDC_GATE_COUNTER 550

`define MODE_PREDICT 	2'b00
`define MODE_TRAIN		2'b01
`define MODE_UPDATE 	2'b11

`define ceilLog2(x) ( \
(x) > 2**30 ? 31 : \
(x) > 2**29 ? 30 : \
(x) > 2**28 ? 29 : \
(x) > 2**27 ? 28 : \
(x) > 2**26 ? 27 : \
(x) > 2**25 ? 26 : \
(x) > 2**24 ? 25 : \
(x) > 2**23 ? 24 : \
(x) > 2**22 ? 23 : \
(x) > 2**21 ? 22 : \
(x) > 2**20 ? 21 : \
(x) > 2**19 ? 20 : \
(x) > 2**18 ? 19 : \
(x) > 2**17 ? 18 : \
(x) > 2**16 ? 17 : \
(x) > 2**15 ? 16 : \
(x) > 2**14 ? 15 : \
(x) > 2**13 ? 14 : \
(x) > 2**12 ? 13 : \
(x) > 2**11 ? 12 : \
(x) > 2**10 ? 11 : \
(x) > 2**9 ? 10 : \
(x) > 2**8 ? 9 : \
(x) > 2**7 ? 8 : \
(x) > 2**6 ? 7 : \
(x) > 2**5 ? 6 : \
(x) > 2**4 ? 5 : \
(x) > 2**3 ? 4 : \
(x) > 2**2 ? 3 : \
(x) > 2**1 ? 2 : \
(x) > 2**0 ? 1 : 0)

`define CELLULAR_AUTOMATON_SEED `HV_DIMENSION'b0001100000000101110111110110000011111100010100111111000000011110100100110110111011110111010101000110101101110110010111111101111100110000011101100111110010000010111111100010001011111100100100000100110011011111000011111000001110000110000010000101000100101111011100110001101100000111010011110100111110001101111010100100000110110111111000111111010010110010011000111111101011110101101001010110110110010111110100100110100010111101000000110011111101000010100011100110100011100110011100011110001110111000000110110100001100011101111100000101110001110001010010100111010101101011110010011011101101010101100111110000101100101001110010011001001010011111101000011010100011011111101011000100000111111010010011111001110110000010110011111110110010011001000100101011100001001101111001011110101111110101111000001111010010001000000100101111011110110101011000111001111111011101100100101010011010001100111100011010010101101101001100101100010011100110111010000011111101001101111111001100001111110101110000111101100110111111

`define BUNDLE_CONNECTIVITY_MATRIX_WIDTH 80000

`define BUNDLE_CONNECTIVITY_MATRIX `BUNDLE_CONNECTIVITY_MATRIX_WIDTH'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111010011110110101100100110100100110110001100111100011111100110100000100001010101100110111111100000011001100001010101010010000000000111000000110010110010001010110011100011000111100110100010101011110100111111111110100110000001101101110010011010000001101010100100001100101100001011100011110010111000111111101111001101001100100100011110110011111000001100101000010001111101110101110001110000001000001101110101011011110101011100111001010010111110100000110011111010011110010010011010111001101101111010100001111001101100000101101001000110010000000000101001111010110001110111000110000000011011110011010010000011111110101000000111010111101011110001100101100111000111000100111000111001001010101000001011111000000011101010001000111001101111000110000111001000010110001000010101000111001000011101101110111011111110001111101101000011100111011100010011100011101001001111001001000001111110111001111000111110111011000110001000111101100001111101100011111100100000010010110110000010001101110001010001101000111111000010000010010111000111000000010010000000111011010001001001000001101000010000001000000110100101100011110011011000000000110010001010001011001110000010000101100100011001101000011000011011100010001100100000110001000100000101000000000100001011100010000000000100000011100000010000110100010011001000000000000001101000011111011000100010101001111110001000100001001011100000010001011110000001111100010000001000001111110100010001010011010010001011010100001010100001000101000101100000100100100000001000010101000000100000010000101101000000000010000101001110000011110010000101110100110000101110011100001010010101110011000100101000101001010100011000000000100001010000001010010110001101010110011011000100011000110101100101101000100000100010100010000100001001110100010000010000110001000000101000000110000010011010010100000100011100001001010001001000011010000001001001010001010000010100010000000000100110001000010110000001000100001001010000000000000110100001001000110011110001000000000100100010001101001001110010001000010000101110100010000110100010000000000000000000000010111000000010101111001011000000000100100000010000000110101000010000100100000000011000001000000000010000111100000001100101000100000000000010000100000000010000000010000000010101000000000100001000001100010010000000110101000100100001000001000100000000110101001001010100011011001000000010000000011000001000110101100000000000100100110001010001000000000001100000000100100010000010010011010100100000000100000100000000000001010101100000000010101000000010000100110000000000100101000100010000101000001101110000010100001000101000100000000000000100000000000101100000010001001001000000101100000000000000100000001001110010010111110010010010000010111111100000010010000100010100010001000001011010000000000000000000010001000000000000001000001000010000001100000010100010001010000000010111000111010000000100000110001000000010000000010010011100100001101100101000000001000000001010000010001000000000101010110100000000100100100001000000100001001000000000001111110001001000110001000000000001001010001000000000001000000000000010000100000001110000000000001101101100100000100100010000000000000000000001000000001100001010000001000000001001001000100000000000001000000100100001000010000000100010001001001100000010010010000000110000000000010001000000000000100100001001000010110010000001000000000010001100000000000101011110001010001011000010000000010001100100000000001000000000000100000000000000000000000000010000000000001000011000001000000010001000000000001011010100001001001000000000010100010000100001010000001000000001101001001000000000000000000011000001000010000001100000000000100000100000011100000000010001000000000000010001010000000001011010010001000101101101000000000000110001000000101010000100000000111000100000000000001000000000000110000000000100010000001000000000000000001001001100000010000100010010000001000000010000100000000001000011001010001000000010000000100000011110000010000000000001001010100000100100000000110000100000110100000010000001000100001111000001000001110000000000000001000000000111110110000000010000010000000000000100001000000100001000001000001000000000000100000000000101000010000001000000000010000000000000000010010110011100000101000000000000010100000000010000100100010100100100000000100101000001001000000001000101010000000000000000110000000001000000000000000000100001000000000100000010011010010001001001001000000000000001111000000001100010000100100000000100000000010101000000000010101010001000000000000000000000000000000101000010000001000001001010000000001011001000100000000000100010010000000000100000011000000000000000000000010100111000000000010001000000001000000000011100000001000100000101000001010000001000000001111010010000000000000000000010001001010000000000010000000000000000000001000000001010001000000000100010010001000000000000000100000010000000100001101000010100001010000000001000000100000000000011000000000001000000000000000100000000000000100000000000000000001001100000000110000000000000000010000011000000001100000000000000000000000100100001011000010000011100010000010000010110000000010000001000000001000001001000000100001000000000000010000001000001000000000000000010000000000000000100001000010100000000100000000000000000000000000000000000001000000000000000000000000000000000000101000000000000001000000100000001000110000010000000000000000010000000000001010000000000000000011100000010000100000001000011010000000100000000101000000001000000000000010001000000001010100000000100000000001010001000000010000000000001000001000000000000000010000000101010000000100000001000000011000000000101110000100000000000100000000010000001000000100000000101000000000000000001000000000000000000000000001100000010100001000000001000000000000000010100100000000000111011100000001000000000010000000100000101000000110000000100000000000000000000100010000010000001100001001001001000000010000001000000010010000000000000100000000000000000000000000110000100000000100000101010111001000000000001000000001010000000000000000001000010000000000000101000001001000001000001000000000000000000100100101000100010000001000010000000000010000001000000001000000000000010000000100000000100000000000000000000000001000000100010000000000000001000000101000010000100000000000000000011000001010000100000000000010010101000010000000000100000000110000000000000001000010000000000000001000000000000000000000000000101001100000000000000001100000000000001110001000000001000101000011100000100000000000000000001000000000010000000000000101000000100000000000010000000000001000001001000000000101000001000010100000000000000000000000100000000100010000000000000100000100000000000011000000000100010000011000000000010000000000000011000000000000101000001000000000000000000100001000000010001010010000000100011000000000000000000000000100000000100000000010010000000101001000000001000001000000000000010000001100000000000000000010000001000000001000010000001000010000000000001000000110000000010000000000000000000010000001000000001000000000000000000000000000000000001000000000110000000000001100000000000000000000000000000000010010000000000000010000000010000010000000001000000000000000101010000100000001000000000000000000000001000000000000001000100001000000000000100000000000000100000000000001000100000001000100000000000000000000001100000000000000000000000000000100001000000110010000000000000100000100000000000000000000010000000000010011110000000000000110101000000000000000000000000001010000000000100001000010000000000000100001000000000000000000000100000010011000000100000000000000000010000000000000000000010000010000000000011000000000000010100000000000000011110000000000000000000000000010000000000000000000000000000001000000000000100001000000000000000001001100000001000000100010000010000000000000000000000000000010010000000000010000001001000000000000001000010000000000000000000000000101000000000000000000000000000000000000000000000110000000001000000000000000000000000000000010000000101001011000101010001010010000010000000100000000001000001000100000000000000000000001001001100000000000000000000000000000100101000000100000000011000000000000000000010000010000100000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000001001000110000000100000110100001000000000010001000000000101000000100001100000000000000000000000001000000000010000000000110001000000010000000000001101000000000100010001000100011000000000000001000000010000010000000000001000000000000000111000000001010000001010001000000000000001110000100000000000100000010000000000000000000000000000000000000000011000000000001100000000000001000000010000000100000000000000000000000010001000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000100001000000000000000000000000000001000000000000001000000000001000000000000100000000010000000000000000000100000000100000000100001000000000010000001000000010000000000010000100000000000000000000100000000000000010100010000000100000000100010000000000001000000000001000000000000001101000000100000000000000001000000010000100000000000000000000000000000000000001000000000000000000000100000000000001000000000000100001000010000000001000010000100000000000000001000000000000000000000010000100000000100000000001000010001000000000000000100000010001000000000010000000000000000001000000001000000000000000100001100000010000000000000001001000000000000001000000000000010000000000000000000000000000000000100000001000000000000000000000000001100000000000000000000000000000000100000110001010001000100000010000000000000000000000000000010000001110010000000000000000000000000000000000010100010000000000000000000000000000100001000000100100000000000000000001000000010010000100000000000100001000000100000000110000000000001000000000001000000001000000001000000001000000000000000100000000000100000000010000000000000000000000000000000000001000010000010000010000000000000000000000110000000000000000000000000100000000000000000000001000000000000000000000001011000000000000000000010000000000000000000010000001000000000000100001000000000000000001000000000000100000000000000000011100000000000000000101000000000100000010000000000000000010100000000011000000000000000000000000000000000000000000100000000000000000100000001100000000000000000000000000101000000000000000100001000000100000000000000000000000000010000000000000000000000000000000000000001000100001000001100000000000000000000000000000001000100001000000000000010000000000000000000000000000100000000000000001010000010010000000000000000000000000000000010000000000000000010000000001000100000000000000000000100000000100000000000000000000000000100010100000000010000010000001001010000000000000000000000000100000000000000000000000000100000000000000000100100000000000000000100000000101000000000000000000000000000001100000000001010100000100000000000000000101100010000000000000000000000010000000000000000000000000000010000100000000000000000000000000000000000000000000000000000001000000000000000000001000000000000000100000000000000000000000000001000100000010000001000000000001000000000001000001000000001000000000000101000000001000010000000000000000001001001000000000001010000000000000000000000000000011000000100000000000000001000010000000000000000000000000010001101000000000000000000000000000100000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000100000110010000000001000000000000000001000001000000001000001000100000000000000000110000000000000000000000000100000000000000000000000001110000000000000000011000011000000000000000000000000000000000000001000000000000000100000000000000000000100000000000000000000000010000000000000000100000000000000000000010000010000011000000100000000000000000000000000000000000001000000000000000000000001000000000001000000000000000000011101000000000000001000000010000000010000010000000000000000000011000000000001000000000000000000100000100000100000000000000000100000000000000000000010000100000010000010000000000000001000000000000100000001000000000000000000000000000000000000000000000000000000000000000001000110000000000000100000000000000000000000000001000000000000000010000000100000000001000000000000100000000000000000000001010000000000100000000010000000000001000000010000000000000100000001001000000000000000000000000100000000000000000011000000000000011000000000000000001000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000101000000000000000010000000000000000000000000000000110000000001000000100000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000100000100000000000000000000000010000000000001010101000000001000000000000001000010000000000000000000000000000100000100000000001101000000000001000000000000100000000000010000000000000000100000000001001000000001010010000010000000000010000000000000001000000100100000000010000000000000000000000001000000000001000001000001000000000000000000010000000000000000000000000000000000000000000010000000000000000000100100000000000000000000000000000010000100000100000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000010000000000000000000000000000000010000000000100000000000000000000000000000000000100000100100000000000001001001000000000000000000000000000000000000000000000000000001000000011000000001001010000000000100000000000000000000000000000000000010000010000000100000000001000100000000000000010100000000000010000000000000001000000000000000000000101000010100000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000100000100000000000001000000000001000000000000010100000000000000000000000001000000000000000000100000000000000000000000000000000000000001000000000000000010000000000000000000000010000000000000000000000000000001000000000000000000000000011000100000001000000000000001010000010000000010000000000010000000001000000000100000100000100000000000010000000000000000000000000000000000000000001000000000000000000000000000001000000000010000000000000000011000000000000000000000000000000000000100000001010000000000000001000010000000000000000000000000000000000000000000010000000000000000000000000100000000000100000000000000000000001000000000000000000000000000100000000001100000000100000000000000000000000000000000100000100000000000000000000001000000000000000000010000000000000000001000000000000000001000000000000000000000000000000000000000000000001000000001000100000100000000000000000000000100000000000000000000000011000001100000010000000010000100000000000000100000000000000000000000000000000000000000000000000000010000100000000000000000011000010000000000000000010000001000000001000100000000000000000000001000000000000000000000000000000000001000000000000000000000000100000000000000000010000010001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000110000000111000100000001000010000000000000000000000000000000010000000000000000000000000000010000000000000000000000010000000000100000000000000000001000010000000000000000000000010000000000000000000000000000010000000010000000000000000000000000000000000110000100000000000000000000000000100000000010000001000000000000000010100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000100000000000000000000000000010000100000000101001000000000001000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010100000010000000010100000000000000100000000000010100000000000010000000000000000000000000000000000000000000001000000000100010000000001000000010000000010000000001000000000000000000001010000000000000000000000000000000000000000000001000000000000000010000110000000000100000100000000000000011000010000000000000000000000001000000000000000000000000000000001000000000000000000000010000010101000000001000000000000000000000000000000000100000000001010000000000000000000000000000000010100000000000000000100000000000000100000010000001010000000000000100000000000000100000000000100000000100001000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000010000000000000000000000100000000000010100000000000010000000000001001000100000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000100000000000000000000000001000000000001000000000000100000000000000000000000000000000010000000000000000000000010000000010000000000000001000000000000001000000010000000001000000000000000000000000000000010000000010000000000000000000000000100000000100000000000000000000000000000000000000000000000000100000100001000101000000010000000000000000000000000000000000000000000000001000000000000000000000000000000010000000001000000100000000000000000000000010000000000000000000000000000000000000000000000000000001010000000000000000000000000000000010000000000000110000000000010000000000001000000001000000000000001100000000000000100000000000100000001000000000000000000000000000000000000000000000000000010000000010010000000000000001010000000000000000000000000000000000000000100000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000010101000110000000000000000000100000100000000000000000000000000000000001000000000000000000000000000001000000000000010000000000000000000000010000000000000000000000000000000000000100000000000000000010000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000110000000010000010000010000000000000000000010000000000000000000000000000000000000000000001001000000000000000000000000000000100000000010000000000000000000001001000000010000000000000000000001000000000000000000000000000001010000000000000000000000000000000100000000001000000000000000000001000000000000000000100000000000010000000000000000000000000000000000000000001000000001000000000001100000000000000000000010000001000000000000110000000010000100100000000000000000000000000000000000000000000010000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000100100100000100000000000000000010000000000000000000010000010000000000000000000000000000001000000000000110000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000001000000000000000000000000010000100000000000000000000000000000000010000000000000000000100000000000100010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000010000100000000000000000001010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000001000000000000000100000000000000000000000000000000000000000001000100000000100000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000110000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001001100000000000000110000000000100010000000000000000000000000000010001100000000000000000000000000000000000000000000000000000000000001000000000000000000001000000010000000000000000000000000000010000000000000000000000000000100010100000000000001000000000000000000000000000000000000000000111000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000001000000000001100000000000000000010000000000000000000000000000010000000010000000000000000100000000000000000000000000000000000000000010010000000000000000000000000000000000000000001000000000000100001000000000000000100000000000000001000000000000000000000000000000000000010000000000000000000000000001000000000000000010000000000000000001000000000000000000000000000000000000000000000100000000000001000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000100000000000000000000000010000000000000000100000000000000000000000000000000001000000100000000100000010000000010000000000000000000100000000000000000000001000000001110000000010000000000000001100000000000000000000000000000000000000000000001000000001000001000100000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000101000000000000100000000000000100000000000000000000000000000000000000000000000000000000000001101000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000001000010000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000100000000000000000000000000000000010000000000000000000000100000000100000010010000000000000000000000000000000000000000001001000000000000000000000000001000000000000000000000010000000000010000000000000000000000000000000000000011000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000100001000000010000000000000000000000100000000000000000000000000000000000000000101000000000001000000000000100000000000000000000000000000000000000000001000001000100000000000000010000000000000000000000000000100000000100000000000000000000000000000000000010000000000000000000001000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000001000000000011000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000001011000000000010000000001000000000000010000001000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000011000000000000000000000100000000000000000000000000000000000000001000000000100000000000000001000000101000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000011000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000010000000000000000000000000000000000100000000100010000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000010000001000000000000000100000000000001100000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000001010000000000000000000000000000000001000000001000000000000000001000000010001000000000000000000000000000000000000000000000000000000000110000000000100000000000001000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000011000000000000000000000010000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000110010000000000000000000000000000000000000010000000000000000000000001000000001000000000000000000000000000000010000000000000000000000000000000000001001000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000010000000000000000000001000000100000001000010000000000000000001000000000000000000010000000000000000000000000000000000000010000000000001000000000000000000000000000000000000000000010000000000000100000000100000000000000000010001000000100000000000000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000010000100000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000001000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000001000000000000000000000000000000100000000000101000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000100000010000000000100000000000010000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000001001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000011000000000000001000001000000100000000010000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000110100000000000001000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000100000000000000000000100000000000000000000000000000000000000100100000000000000000001000000000000000000000000000000000100000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000010000000000010000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000010000000000000000000100000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000001000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000100000101000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100000000000000001000000000000000000000000000000000000010010000000000000000000100000000100000000000000000000000000010000000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010011000000000000000000000000000100000000001000000000100000010000000000000000000000100000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000010101000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000100001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000001000000000000000000000000000000100000000001000000010000000000000000000000000000000000000000000010000000000000000000010000000001000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000010000010000100000000000000000000000000000000000000100000000000000000000001000100000000000000000000100000000000000000000100000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000100010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000010100000000000000000000000010001000000000001000000000100000000000000000000000000000000000100000000000000000000000000100001000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000010000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000001001010000000000000000000000000000000101000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000001000000000000000000000010000000000000000000000000010001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000001000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000010000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000100000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000010000000100000100000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100010100000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000100000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000001000000000000000001100000000000000000000000000000000100001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000000000100000100000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000100000010000000001000000000000000000000000000000000000000000000000000000000000000000000110000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000001000000010000000001000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000010000000000000000000000000000001000010000000000000000000000000000000000000000100000000000001000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000010000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000010000000010000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000001000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000100000000000000000010010000000000000000000000000000000000000000100000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000010000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000100000000000100000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000001000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000100000000000000000000000000000001000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000100000000000000000000000010000001000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000011000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000001000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000010001000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000100000000000010000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000100001000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000001000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000001000000000000000000000010000000000000000000000001000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000001000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000100000000100000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000010000000000000100000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000110000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000110000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000000000000000000000000000000000000000100000001001000000100010000100000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000001000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000100000000100000000000000000010000000000000100100000000000000000000000000000000001010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010011000000001010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000010000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000010000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000001000000000001000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000001000000100000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000100000000010000000001000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000100000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000001000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000001000000000000000100000000000000000010000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000100000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000010000000000010000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000100000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000010001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000010000000000000000000000010001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001010000000000000000000000000000000000000010000000000000000000000000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000001000000000000000000000000000000000000110000000000000000000100000000000000000000000000000000000000000000000011000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000010000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000100000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000001000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000100010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001010000000000000000000000000010000000000000000000000000000000010000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000100000010000000000000000000000000000000000000000000000000001000100000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010001000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000

`define MERGE_BITS `HV_DIMENSION'b1111101100001010001101000111001110100111111010110010010010010000100111111000111010011100010110101001010100010101001001000100010011000100001011111100010000010011001100010101011010100011010010011010010100001001110101011100111001101111100101000100000100100001000011010000011010000111000011000111101101100010011100111001000111001101001000000100010111000111111010001001011000001101110001001111101010001100010111001111111011111000101100000010000100100001001010111110111001010011000111100101100011010101100110001000001011100110001101101000000111100100111100000001010000110110111011111010001111100101101101110110011010001100011010101001111011011001000011111101011001111001100001101101010100100110100111100111101110101011101101010110100111010110000100000000010010000000000001111011111010000110011110110111011100111100000111000110000100110111000100001111111011110101111100110100110111010111111111010101111001100100101110101111110111110100001000110001110010100010011000000110011110001110101111100111100011011101

`endif