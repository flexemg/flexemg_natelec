//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Sat Feb 04 07:43:01 2017
// Version: v11.7 SP3 11.7.3.8
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// mux_2x_2_1
module mux_2x_2_1(
    // Inputs
    A0,
    A1,
    B0,
    B1,
    SEL,
    // Outputs
    Y0,
    Y1
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  A0;
input  A1;
input  B0;
input  B1;
input  SEL;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output Y0;
output Y1;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   A0;
wire   A1;
wire   B0;
wire   B1;
wire   SEL;
wire   Y0_net_0;
wire   Y1_net_0;
wire   Y0_net_1;
wire   Y1_net_1;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign Y0_net_1 = Y0_net_0;
assign Y0       = Y0_net_1;
assign Y1_net_1 = Y1_net_0;
assign Y1       = Y1_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------MX2
MX2 MX2_0(
        // Inputs
        .A ( A0 ),
        .B ( B0 ),
        .S ( SEL ),
        // Outputs
        .Y ( Y0_net_0 ) 
        );

//--------MX2
MX2 MX2_1(
        // Inputs
        .A ( A1 ),
        .B ( B1 ),
        .S ( SEL ),
        // Outputs
        .Y ( Y1_net_0 ) 
        );


endmodule
